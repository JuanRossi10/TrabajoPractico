library verilog;
use verilog.vl_types.all;
entity Sec_LED_vlg_vec_tst is
end Sec_LED_vlg_vec_tst;
