library verilog;
use verilog.vl_types.all;
entity EjercicioLED_vlg_vec_tst is
end EjercicioLED_vlg_vec_tst;
