library verilog;
use verilog.vl_types.all;
entity Block1_vlg_check_tst is
    port(
        Q               : in     vl_logic;
        Q35             : in     vl_logic;
        Q36             : in     vl_logic;
        Q37             : in     vl_logic;
        Q38             : in     vl_logic;
        Q39             : in     vl_logic;
        Q40             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Block1_vlg_check_tst;
