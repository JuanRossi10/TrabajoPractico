library verilog;
use verilog.vl_types.all;
entity Block1 is
    port(
        clock           : in     vl_logic;
        D               : in     vl_logic;
        D41             : in     vl_logic;
        D42             : in     vl_logic;
        D43             : in     vl_logic;
        D44             : in     vl_logic;
        D45             : in     vl_logic;
        D46             : in     vl_logic;
        D47             : in     vl_logic;
        D48             : in     vl_logic;
        Q               : out    vl_logic;
        Q35             : out    vl_logic;
        Q36             : out    vl_logic;
        Q37             : out    vl_logic;
        Q38             : out    vl_logic;
        Q39             : out    vl_logic;
        Q40             : out    vl_logic
    );
end Block1;
