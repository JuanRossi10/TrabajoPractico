library verilog;
use verilog.vl_types.all;
entity Sec_LED_vlg_check_tst is
    port(
        z1              : in     vl_logic;
        z2              : in     vl_logic;
        z3              : in     vl_logic;
        z4              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Sec_LED_vlg_check_tst;
